module memory
#(parameter Data_width = 16, Addr_width = 12)
(
input clk,we,
input [Addr_width-1:0] addr,
input [Data_width-1:0] din,
output reg [Data_width-1:0] dout);

reg [Data_width-1:0] ram [2**Addr_width-1:0];

initial begin
	$readmemb("D:\\Work_Parent\\Octacore Processor\\11-Input_handler\\Memory_file.txt",ram);
end

/*
initial 
begin
//instructions
ram[0] = 16'b1110000000000000;
ram[1] = 16'b1110000000000000;
ram[2] = 16'b1110000000000000;
ram[3] = 16'b1000000000000000;
ram[4] = 16'b0000111110100000;
ram[5] = 16'b0000111110100001;
ram[6] = 16'b0000111110100010;
ram[7] = 16'b0000111110100011;
ram[8] = 16'b0001111110100101;
ram[9] = 16'b0110000000000000;
ram[10] = 16'b0001111110100000;
ram[11] = 16'b1011000000000000;
ram[12] = 16'b0110000000000000;
ram[13] = 16'b0001111110100010;
ram[14] = 16'b1001000000000000;
ram[15] = 16'b0110000000000000;
ram[16] = 16'b0001101110111000;
ram[17] = 16'b1001000000000000;
ram[18] = 16'b0011000000000000;
ram[19] = 16'b0111000000000000;
ram[20] = 16'b0100000000000000;
ram[21] = 16'b0001111110100010;
ram[22] = 16'b0110000000000000;
ram[23] = 16'b0001111110100110;
ram[24] = 16'b1011000000000000;
ram[25] = 16'b0110000000000000;
ram[26] = 16'b0001111110100001;
ram[27] = 16'b1001000000000000;
ram[28] = 16'b0110000000000000;
ram[29] = 16'b0001101110111001;
ram[30] = 16'b1001000000000000;
ram[31] = 16'b0011000000000000;
ram[32] = 16'b0101000000000000;
ram[33] = 16'b1011000000000000;
ram[34] = 16'b0100000000000000;
ram[35] = 16'b0001111110100011;
ram[36] = 16'b0110000000000000;
ram[37] = 16'b0001101110111010;
ram[38] = 16'b1001000000000000;
ram[39] = 16'b0011000000000000;
ram[40] = 16'b0101000000000000;
ram[41] = 16'b1001000000000000;
ram[42] = 16'b0100000000000000;
ram[43] = 16'b0001111110100011;
ram[44] = 16'b0110000000000000;
ram[45] = 16'b0001101110111010;
ram[46] = 16'b1001000000000000;
ram[47] = 16'b0110000000000000;
ram[48] = 16'b0101000000000000;
ram[49] = 16'b0010000000000000;
ram[50] = 16'b0001111110100010;
ram[51] = 16'b1100000000000000;
ram[52] = 16'b0000111110100010;
ram[53] = 16'b0110000000000000;
ram[54] = 16'b0001111110100101;
ram[55] = 16'b1010000000000000;
ram[56] = 16'b1101000000001000;
ram[57] = 16'b0000111110100010;
ram[58] = 16'b0001111110100011;
ram[59] = 16'b1100000000000000;
ram[60] = 16'b0000111110100011;
ram[61] = 16'b0001111110100001;
ram[62] = 16'b1100000000000000;
ram[63] = 16'b0000111110100001;
ram[64] = 16'b0110000000000000;
ram[65] = 16'b0001111110100110;
ram[66] = 16'b1010000000000000;
ram[67] = 16'b1101000000001000;
ram[68] = 16'b0000111110100001;
//ram[69] = 16'b0000111110100010;
ram[69] = 16'b0001111110100000;
ram[70] = 16'b1100000000000000;
ram[71] = 16'b0000111110100000;
ram[72] = 16'b0110000000000000;
ram[73] = 16'b0001111110100100;
ram[74] = 16'b1010000000000000;
ram[75] = 16'b1101000000001000;
ram[76] = 16'b1110000000000000;
ram[77] = 16'b1111000000000000;

//m
ram[4004] = 3;
//q
ram[4005] = 3;
//n
ram[4006] = 3;
//baseA
ram[3000] = 3800;
//baseB
ram[3001] = 3850;
//baseC
ram[3002] = 3900;
//A
ram[3800] = 1;
ram[3801] = 2;
ram[3802] = 3;
ram[3803] = 4;
ram[3804] = 5;
ram[3805] = 6;
ram[3806] = 7;
ram[3807] = 8;
ram[3808] = 9;
//B
ram[3850] = 2;
ram[3851] = 3;
ram[3852] = 5;
ram[3853] = 7;
ram[3854] = 11;
ram[3855] = 13;
ram[3856] = 17;
ram[3857] = 19;
ram[3858] = 23;


//C
ram[3900] = 0;
ram[3901] = 0;
ram[3902] = 0;
ram[3903] = 0;
ram[3904] = 0;
ram[3905] = 0;
ram[3906] = 0;
ram[3907] = 0;
ram[3908] = 0;
ram[3909] = 0;
ram[3910] = 0;
ram[3911] = 0;

end
*/

always@(posedge clk)
begin
if(we)
begin
	ram[addr]<=din;
end else begin
	dout<=ram[addr];
end
end

endmodule